library IEEE;
use IEEE.std_logic_1164.all;
library LIB_AES;
use LIB_AES.Crypt_Pack.all;

entity SBox is
    port (
        SBox_i : in bit8;
        SBox_o : out bit8);
end entity;

architecture SBox_arch of SBox is

begin
P1:process (SBox_i)
begin
    ---les colonnes de Sbox
    case SBox_i is
        when X"00" => SBox_o <= X"63";
        when X"10" => SBox_o <= X"ca";
        when X"20" => SBox_o <= X"b7";
        when X"30" => SBox_o <= X"04";
        when X"40" => SBox_o <= X"09";
        when X"50" => SBox_o <= X"53";
        when X"60" => SBox_o <= X"d0";
        when X"70" => SBox_o <= X"51";
        when X"80" => SBox_o <= X"cd";
        when X"90" => SBox_o <= X"60";
        when X"a0" => SBox_o <= X"e0";
        when X"b0" => SBox_o <= X"e7";
        when X"c0" => SBox_o <= X"ba";
        when X"d0" => SBox_o <= X"70";
        when X"e0" => SBox_o <= X"e1";
        when X"f0" => SBox_o <= X"8c";

        when X"01" => SBox_o <= X"7c";
        when X"11" => SBox_o <= X"82";
        when X"21" => SBox_o <= X"fd";
        when X"31" => SBox_o <= X"c7";
        when X"41" => SBox_o <= X"83";
        when X"51" => SBox_o <= X"d1";
        when X"61" => SBox_o <= X"ef";
        when X"71" => SBox_o <= X"a3";
        when X"81" => SBox_o <= X"0c";
        when X"91" => SBox_o <= X"81";
        when X"a1" => SBox_o <= X"32";
        when X"b1" => SBox_o <= X"c8";
        when X"c1" => SBox_o <= X"78";
        when X"d1" => SBox_o <= X"3e";
        when X"e1" => SBox_o <= X"f8";
        when X"f1" => SBox_o <= X"a1";

        when X"02" => SBox_o <= X"77";
        when X"12" => SBox_o <= X"c9";
        when X"22" => SBox_o <= X"93";
        when X"32" => SBox_o <= X"23";
        when X"42" => SBox_o <= X"2c";
        when X"52" => SBox_o <= X"00";
        when X"62" => SBox_o <= X"aa";
        when X"72" => SBox_o <= X"40";
        when X"82" => SBox_o <= X"13";
        when X"92" => SBox_o <= X"4f";
        when X"a2" => SBox_o <= X"3a";
        when X"b2" => SBox_o <= X"37";
        when X"c2" => SBox_o <= X"25";
        when X"d2" => SBox_o <= X"b5";
        when X"e2" => SBox_o <= X"98";
        when X"f2" => SBox_o <= X"89";

        when X"03" => SBox_o <= X"7b";
        when X"13" => SBox_o <= X"7d";
        when X"23" => SBox_o <= X"26";
        when X"33" => SBox_o <= X"c3";
        when X"43" => SBox_o <= X"1a";
        when X"53" => SBox_o <= X"ed";
        when X"63" => SBox_o <= X"fb";
        when X"73" => SBox_o <= X"8f";
        when X"83" => SBox_o <= X"ec";
        when X"93" => SBox_o <= X"dc";
        when X"a3" => SBox_o <= X"0a";
        when X"b3" => SBox_o <= X"6d";
        when X"c3" => SBox_o <= X"2e";
        when X"d3" => SBox_o <= X"66";
        when X"e3" => SBox_o <= X"11";
        when X"f3" => SBox_o <= X"0d";

        when X"04" => SBox_o <= X"f2";
        when X"14" => SBox_o <= X"fa";
        when X"24" => SBox_o <= X"36";
        when X"34" => SBox_o <= X"18";
        when X"44" => SBox_o <= X"1b";
        when X"54" => SBox_o <= X"20";
        when X"64" => SBox_o <= X"43";
        when X"74" => SBox_o <= X"92";
        when X"84" => SBox_o <= X"5f";
        when X"94" => SBox_o <= X"22";
        when X"a4" => SBox_o <= X"49";
        when X"b4" => SBox_o <= X"8d";
        when X"c4" => SBox_o <= X"1c";
        when X"d4" => SBox_o <= X"84";
        when X"e4" => SBox_o <= X"69";
        when X"f4" => SBox_o <= X"bf";

        when X"05" => SBox_o <= X"6b";
        when X"15" => SBox_o <= X"59";
        when X"25" => SBox_o <= X"3f";
        when X"35" => SBox_o <= X"96";
        when X"45" => SBox_o <= X"6e";
        when X"55" => SBox_o <= X"fc";
        when X"65" => SBox_o <= X"4d";
        when X"75" => SBox_o <= X"9d";
        when X"85" => SBox_o <= X"97";
        when X"95" => SBox_o <= X"2a";
        when X"a5" => SBox_o <= X"06";
        when X"b5" => SBox_o <= X"d5";
        when X"c5" => SBox_o <= X"a6";
        when X"d5" => SBox_o <= X"03";
        when X"e5" => SBox_o <= X"d9";
        when X"f5" => SBox_o <= X"e6";
        
        when X"06" => SBox_o <= X"6f";
        when X"16" => SBox_o <= X"47";
        when X"26" => SBox_o <= X"f7";
        when X"36" => SBox_o <= X"05";
        when X"46" => SBox_o <= X"5a";
        when X"56" => SBox_o <= X"b1";
        when X"66" => SBox_o <= X"33";
        when X"76" => SBox_o <= X"38";
        when X"86" => SBox_o <= X"44";
        when X"96" => SBox_o <= X"90";
        when X"a6" => SBox_o <= X"24";
        when X"b6" => SBox_o <= X"4e";
        when X"c6" => SBox_o <= X"b4";
        when X"d6" => SBox_o <= X"f6";
        when X"e6" => SBox_o <= X"8e";
        when X"f6" => SBox_o <= X"42";
        when X"07" => SBox_o <= X"c5";
        when X"17" => SBox_o <= X"f0";
        when X"27" => SBox_o <= X"cc";
        when X"37" => SBox_o <= X"9a";
        when X"47" => SBox_o <= X"a0";
        when X"57" => SBox_o <= X"5b";
        when X"67" => SBox_o <= X"85";
        when X"77" => SBox_o <= X"f5";
        when X"87" => SBox_o <= X"17";
        when X"97" => SBox_o <= X"88";
        when X"a7" => SBox_o <= X"5c";
        when X"b7" => SBox_o <= X"a9";
        when X"c7" => SBox_o <= X"c6";
        when X"d7" => SBox_o <= X"0e";
        when X"e7" => SBox_o <= X"94";
        when X"f7" => SBox_o <= X"68";
        when X"08" => SBox_o <= X"30";
        when X"18" => SBox_o <= X"ad";
        when X"28" => SBox_o <= X"34";
        when X"38" => SBox_o <= X"07";
        when X"48" => SBox_o <= X"52";
        when X"58" => SBox_o <= X"6a";
        when X"68" => SBox_o <= X"45";
        when X"78" => SBox_o <= X"bc";
        when X"88" => SBox_o <= X"c4";
        when X"98" => SBox_o <= X"46";
        when X"a8" => SBox_o <= X"c2";
        when X"b8" => SBox_o <= X"6c";
        when X"c8" => SBox_o <= X"e8";
        when X"d8" => SBox_o <= X"61";
        when X"e8" => SBox_o <= X"9b";
        when X"f8" => SBox_o <= X"41";
        when X"09" => SBox_o <= X"01";
        when X"19" => SBox_o <= X"d4";
        when X"29" => SBox_o <= X"a5";
        when X"39" => SBox_o <= X"12";
        when X"49" => SBox_o <= X"3b";
        when X"59" => SBox_o <= X"cb";
        when X"69" => SBox_o <= X"f9";
        when X"79" => SBox_o <= X"b6";
        when X"89" => SBox_o <= X"a7";
        when X"99" => SBox_o <= X"ee";
        when X"a9" => SBox_o <= X"d3";
        when X"b9" => SBox_o <= X"56";
        when X"c9" => SBox_o <= X"dd";
        when X"d9" => SBox_o <= X"35";
        when X"e9" => SBox_o <= X"1e";
        when X"f9" => SBox_o <= X"99";
        when X"0a" => SBox_o <= X"67";
        when X"1a" => SBox_o <= X"a2";
        when X"2a" => SBox_o <= X"e5";
        when X"3a" => SBox_o <= X"80";
        when X"4a" => SBox_o <= X"d6";
        when X"5a" => SBox_o <= X"be";
        when X"6a" => SBox_o <= X"02";
        when X"7a" => SBox_o <= X"da";
        when X"8a" => SBox_o <= X"7e";
        when X"9a" => SBox_o <= X"b8";
        when X"aa" => SBox_o <= X"ac";
        when X"ba" => SBox_o <= X"f4";
        when X"ca" => SBox_o <= X"74";
        when X"da" => SBox_o <= X"57";
        when X"ea" => SBox_o <= X"87";
        when X"fa" => SBox_o <= X"2d";
        when X"0b" => SBox_o <= X"2b";
        when X"1b" => SBox_o <= X"af";
        when X"2b" => SBox_o <= X"f1";
        when X"3b" => SBox_o <= X"e2";
        when X"4b" => SBox_o <= X"b3";
        when X"5b" => SBox_o <= X"39";
        when X"6b" => SBox_o <= X"7f";
        when X"7b" => SBox_o <= X"21";
        when X"8b" => SBox_o <= X"3d";
        when X"9b" => SBox_o <= X"14";
        when X"ab" => SBox_o <= X"62";
        when X"bb" => SBox_o <= X"ea";
        when X"cb" => SBox_o <= X"1f";
        when X"db" => SBox_o <= X"b9";
        when X"eb" => SBox_o <= X"e9";
        when X"fb" => SBox_o <= X"0f";
        when X"0c" => SBox_o <= X"fe";
        when X"1c" => SBox_o <= X"9c";
        when X"2c" => SBox_o <= X"71";
        when X"3c" => SBox_o <= X"eb";
        when X"4c" => SBox_o <= X"29";
        when X"5c" => SBox_o <= X"4a";
        when X"6c" => SBox_o <= X"50";
        when X"7c" => SBox_o <= X"10";
        when X"8c" => SBox_o <= X"64";
        when X"9c" => SBox_o <= X"de";
        when X"ac" => SBox_o <= X"91";
        when X"bc" => SBox_o <= X"65";
        when X"cc" => SBox_o <= X"4b";
        when X"dc" => SBox_o <= X"86";
        when X"ec" => SBox_o <= X"ce";
        when X"fc" => SBox_o <= X"b0";
        when X"0d" => SBox_o <= X"d7";
        when X"1d" => SBox_o <= X"a4";
        when X"2d" => SBox_o <= X"d8";
        when X"3d" => SBox_o <= X"27";
        when X"4d" => SBox_o <= X"e3";
        when X"5d" => SBox_o <= X"4c";
        when X"6d" => SBox_o <= X"3c";
        when X"7d" => SBox_o <= X"ff";
        when X"8d" => SBox_o <= X"5d";
        when X"9d" => SBox_o <= X"5e";
        when X"ad" => SBox_o <= X"95";
        when X"bd" => SBox_o <= X"7a";
        when X"cd" => SBox_o <= X"bd";
        when X"dd" => SBox_o <= X"c1";
        when X"ed" => SBox_o <= X"55";
        when X"fd" => SBox_o <= X"54";
        when X"0e" => SBox_o <= X"ab";
        when X"1e" => SBox_o <= X"72";
        when X"2e" => SBox_o <= X"31";
        when X"3e" => SBox_o <= X"b2";
        when X"4e" => SBox_o <= X"2f";
        when X"5e" => SBox_o <= X"58";
        when X"6e" => SBox_o <= X"9f";
        when X"7e" => SBox_o <= X"f3";
        when X"8e" => SBox_o <= X"19";
        when X"9e" => SBox_o <= X"0b";
        when X"ae" => SBox_o <= X"e4";
        when X"be" => SBox_o <= X"ae";
        when X"ce" => SBox_o <= X"8b";
        when X"de" => SBox_o <= X"1d";
        when X"ee" => SBox_o <= X"28";
        when X"fe" => SBox_o <= X"bb";
        when X"0f" => SBox_o <= X"76";
        when X"1f" => SBox_o <= X"c0";
        when X"2f" => SBox_o <= X"15";
        when X"3f" => SBox_o <= X"75";
        when X"4f" => SBox_o <= X"84";
        when X"5f" => SBox_o <= X"cf";
        when X"6f" => SBox_o <= X"a8";
        when X"7f" => SBox_o <= X"d2";
        when X"8f" => SBox_o <= X"73";
        when X"9f" => SBox_o <= X"db";
        when X"af" => SBox_o <= X"79";
        when X"bf" => SBox_o <= X"08";
        when X"cf" => SBox_o <= X"8a";
        when X"df" => SBox_o <= X"9e";
        when X"ef" => SBox_o <= X"df";
        when X"ff" => SBox_o <= X"16";        
        when others => SBox_o <= X"63";   
    end case;
end process;

end architecture;